`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:12:50 01/20/2023 
// Design Name: 
// Module Name:    ledrandom 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ledrandom(randominput,ledsout
    );
	 
	 //This module is taking the 4-bit random number
	 //generated by random number generator and lights
	 //the LEDs.For example if the number is 1011 then
	 //first,second and fourth LEDs will light.The reason
	 //i did this module is that i couldn't directly use
	 //the output because in Verilog we can't use 1 input or
	 //output in more than 1 always block in 1 module.
	 input [3:0] randominput;
	 output reg [3:0] ledsout;
	 
	 always @(randominput[0] or randominput[1] or randominput[2] or randominput[3]) begin
	 
	 ledsout = randominput;
	 end
	         

endmodule
